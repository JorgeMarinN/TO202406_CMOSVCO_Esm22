** sch_path: /home/designer/shared/Workshop-CANELOS24/xschem/TB_DCDCBuck_V2.sch
**.subckt TB_DCDCBuck_V2
Vdd Vdd GND 3.3
Vg2 Vg_M2 GND PULSE(0 {VH} {dt} 1n 1n {T*D-2*dt} {T} 0)
Vg1 Vg_M1 GND PULSE(0 {VH} 0 1n 1n {T*D} {T} 0)
XM2 Vc Vg_M2 GND GND sg13_hv_nmos w={w_M2} l={l_M2} ng={ng_M2} m={mult_M2}
XM1 Vc Vg_M1 Vdd Vdd sg13_hv_pmos w={w_M1} l={l_M1} ng={ng_M1} m={mult_M1}
L6 net2 net1 {L} m=1
C1 net1 GND {C} m=1
V_Io net1 Vo 0
.save i(v_io)
V_IL Vc net2 0
.save i(v_il)
R2 Vo GND {R} m=1
**** begin user architecture code


*Parametros
*Filtro
.param L = 1.37u
.param R = 0.9
.param C = 416n





.param temp=27
*.param mult_M1 = 2400
.param mult_M1 = 3600
.param w_M1 =10u
*.param l_M1 = 0.2u ** Posee mayor capacidad de corriente, pero en sub-umbral conduce mucha corriente
.param l_M1 = 0.22u
.param ng_M1 = 1

*.param mult_M2 = 1200
.param mult_M2 = 1800
.param w_M2 =10u
*.param l_M2 =0.25u
.param l_M2 =0.25u
.param ng_M2 =1








.param VH = 3
.param D = 0.42
.param T = 1u
.param dt = 5n
.param temp = 27






.save all
.control
reset
set color0 = white
tran 1n 100u
plot i(V_Io) i(V_IL)
plot v(Vo)
plot v(Vc)
plot v(Vg_M1) v(Vg_M2)
.endc

.end



.lib cornerMOShv.lib mos_tt

**** end user architecture code
**.ends
.GLOBAL GND
.end
